parameter ADDR_WIDTH = 10;//������ ���� �����
parameter DATA_REG_ADDR = 10'd5; //����� �������� ������
parameter CONFIG_REG_ADDR = 10'd6; //����� ����������������� ��������
parameter STATUS_REG_ADDR = 10'd7; //����� ���������� ��������
parameter CONFIG_REG_WIDTH = 8;//������ ����������������� ��������
parameter STATUS_REG_WIDTH = 8;//������ ���������� ��������