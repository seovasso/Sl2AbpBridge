`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12.10.2017 17:57:40
// Design Name: 
// Module Name: ApbSlTb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
parameter clkPeriod=10;//������ �����
parameter clkTimeDiff=3;//�������� �������� �������� ������������ ���� �����
parameter paddrWidth=10;// ������ �������� ���� apb
module Apb2SlTb(

    );

    logic clk; //�������� �������: �����
    logic pclk;// apb
    // ������� ���� apb
    logic                   preset_n;
    logic                   reset_n;
    logic [paddrWidth-1:0]  paddr;
    logic                   pprot;
    logic                   psel2;
    logic                   penable;
    logic                   pwrite;
    logic [31:0]            pwdata;
    logic [31:0]            prdata;
    logic [3:0]             pstrb;
    logic                   pready;
    logic                   pdata;
    logic                   pslverr;
    //����������� ������
         Apb2Sl mod (
          .clk(clk),
          .pclk(pclk),
          .reset_n(reset_n),
          .psel1(psel2),
          .paddr(paddr),
          .pwdata(pwdata),
          .prdata(pwdata),
          .penable(penable),
          .pready(pready),
          .pslverr(pslverr),
          .pstrb(pstrb),
          .preset_n(preset_n)
   );
    
    
    // �������� ���������� ������ � ������
    task writeTransaction;
      input bit [31:0] wrData;
      input bit [paddrWidth-1:0] wrAddr;
      begin 
      #clkPeriod;
        paddr=wrAddr;
        pwrite=1;
        penable=0;
        pstrb=4'b1111;
        pwdata=wrData;
        psel2=1;
      #clkPeriod;
        penable=1;
      #clkPeriod;
      //while(!pready)begin
        psel2=0;
        penable=0;
        pwdata=0;
        paddr=0; 
        pstrb=0;  
        pwrite=0; 
      end
    endtask;
    task readTransaction();
          begin 
          
          end
        endtask;
    
    initial
      begin
       #(clkTimeDiff);
        forever #(clkPeriod/2) clk<=~clk;//������ ����
      end
    initial
      begin
        forever #(clkPeriod/2) pclk<=~pclk;//������ ����
      end
     initial begin
     //�������������
     clk=0;
     pclk=0;
     preset_n=1;
     paddr=0;
     pprot=0;
     psel2=0;
     penable=0;
     pwrite=0;
     pwdata=0;
     pstrb=0;
     #25;
     preset_n=0;
     #15;
     preset_n=1;
     #40
     writeTransaction(10'd2,32'd3156);
     end

endmodule
